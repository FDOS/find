# Translation by Martin Strömberg <ams@ludd.luth.se>.
0.0:Visar alla rader i en fil som innehåller en viss sträng
0.1:Räkna antalet gånger strängen förekommer
0.2:Hantera versaler och gemener som lika
0.3:Numrera de visade raderna med start från 1
0.4:Visa raderna som inte innehåller strängen
1.0:fil
1.1:sträng
2.0:Kan inte öppna filen
2.1:Ingen sådan fil
2.2:Kan inte byta till katalog
